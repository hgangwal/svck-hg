package p1;
  int tt;
endpackage: p1

package p2;
  int i1;
class c;
  rand int t;
  local int lvar_i1;
endclass : c
endpackage: p2
