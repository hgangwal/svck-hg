class c;
  protected int state_snake_name_1;
  rand int camelCaseName2;
  local int PascalCaseName3;
endclass : c

class c2;
  local int state_i1;
  rand int rand_i1;
  local int lvar_i1;
  local int prot_i1;
endclass : c2
