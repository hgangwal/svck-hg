class c;
  protected int state_i1;
  rand int rand_i1;
  local int lvar_i1;
endclass : c

class c2;
  int state_i1;
  rand int rand_i1;
  int lvar_i1;
  int prot_i1;
endclass : c2
