/*
# ----------------------------------------------------
# SPDX-FileCopyrightText: AsFigo Technologies, UK
# SPDX-FileCopyrightText: VerifWorks, India
# SPDX-License-Identifier: MIT
# Author: Saavni Pradhan 
# ----------------------------------------------------
*/
class c;
  mailbox bad_gbx;
  mailbox #(int) good_ibx;
endclass : c
